** Profile: "SCHEMATIC1-PSiNu"  [ C:\Users\Cristi\Desktop\LAB ASCN 1\1-PSpiceFiles\SCHEMATIC1\PSiNu.sim ] 

** Creating circuit file "PSiNu.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\Users\Cristi\Desktop\LAB ASCN 1\1-PSpiceFiles\SCHEMATIC1\PSiNu\PSiNu_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Cristi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
