** Profile: "SCHEMATIC1-DMUX"  [ C:\Users\Cristi\Desktop\LAB ASCN 1\dmux-pspicefiles\schematic1\dmux.sim ] 

** Creating circuit file "DMUX.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\Users\Cristi\Desktop\LAB ASCN 1\dmux-pspicefiles\schematic1\DMUX\DMUX_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Cristi\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 16 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
